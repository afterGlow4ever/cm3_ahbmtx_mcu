//===============================================
//
//	File: fpga_universal_sp_sram_gen.v
//	Author: afterGlow,4ever
//	Date: 05022024
//	Version: v1.0
//
// 	This lib is used to generate fpga universal sram 
// 	including:
// 	1. altera sp ram
// 	2. xilinx sp ram
// 	3. simple sim ram
//
//	The active value of be, we, ce are all high.
//
//===============================================

module fpga_universal_sp_sram_gen
(
	clk,
	rst,
	be,
	we,
	cs,
	addr,
	data,
	q
);

parameter									ADDR_WIDTH = 10;
parameter									DATA_WIDTH = 32;
parameter									BYTE_WIDTH = 8;
parameter									MEM_INITFILE = "none";
parameter									BYTE_RESIDUAL = (DATA_WIDTH%BYTE_WIDTH) ? 1 : 0;
parameter									BYTE_QUOTIENT = (DATA_WIDTH/BYTE_WIDTH) + BYTE_RESIDUAL;
parameter									BYTE_NUMBER = BYTE_QUOTIENT + BYTE_RESIDUAL;
parameter									FULL_DATA_WIDTH = BYTE_NUMBER*BYTE_WIDTH;

input										clk;
input										rst;
input		[BYTE_NUMBER-1:0]				be;
input										we;
input										cs;
input	 	[ADDR_WIDTH-1:0]				addr;
input		[DATA_WIDTH-1:0]				data;
output		[DATA_WIDTH-1:0]				q;

wire		[FULL_DATA_WIDTH-1:0]			real_data;
wire		[FULL_DATA_WIDTH-1:0]			real_q;

assign real_data = {{(FULL_DATA_WIDTH-DATA_WIDTH){1'b0}}, data};
assign q = real_q[DATA_WIDTH-1:0];

//===============================================
// If BYTE_WIDTH is not 8 or 9, this ram will be
// generated by multiple parallel rams.
// If BYTE_WIDTH is 8 or 9, this ram will be
// generated by a single ram.
//===============================================

genvar										i, j;

generate
	if((BYTE_WIDTH!=8)&&(BYTE_WIDTH!=9))
	begin: multi_sp_ram_gen
		for(i=0;i<BYTE_NUMBER;i=i+1)
		begin: sp_ram_gen
`ifdef FPGA_SRAM
`ifdef ALTERA_EP4
			altera_sp_sram_gen
			#(
				.ADDR_WIDTH(ADDR_WIDTH),
				.DATA_WIDTH(BYTE_WIDTH),
				.BYTE_WIDTH(BYTE_WIDTH),
				.MEM_INITFILE(),
				.DEVICE_FAMILY("Cyclone IV E")
			)
			u_sp_sram_gen
			(
				.clk						(clk),
				.rst						(rst),
				.byteena					(1'b1),
				.wren						(we&be[i]&cs),
				.rden						(cs&!we)),//?
				.addr						(addr),
				.data						(real_data[(i+1)*BYTE_WIDTH-1:i*BYTE_WIDTH]),
				.q							(real_q[(i+1)*BYTE_WIDTH-1:i*BYTE_WIDTH])
			);
`elsif ZYNQ_7020
			xilinx_sp_sram_gen
			#(
				.ADDR_WIDTH(ADDR_WIDTH),
				.DATA_WIDTH(BYTE_WIDTH),
				.BYTE_WIDTH(BYTE_WIDTH),
				.MEM_INITFILE(),
				.DEVICE_FAMILY("ZYNQ_7020")
			)
			u_sp_sram_gen
			(
				.clk						(clk),
				.rst						(rst),
				.wea						(we&be[i]),
				.ena						(cs),
				.addr						(addr),
				.data						(real_data[(i+1)*BYTE_WIDTH-1:i*BYTE_WIDTH]),
				.q							(real_q[(i+1)*BYTE_WIDTH-1:i*BYTE_WIDTH])
			);
`else
`endif
`else
			sim_sp_sram_gen
			#(
				.ADDR_WIDTH(ADDR_WIDTH),
				.DATA_WIDTH(BYTE_WIDTH),
				.BYTE_WIDTH(BYTE_WIDTH),
				.MEM_INITFILE()
			)
			u_sp_sram_gen
			(
				.clk						(clk),
				.rst						(rst),
				.wea						(we&be[i]),
				.ena						(cs),
				.addr						(addr),
				.data						(real_data[(i+1)*BYTE_WIDTH-1:i*BYTE_WIDTH]),
				.q							(real_q[(i+1)*BYTE_WIDTH-1:i*BYTE_WIDTH])
			);
`endif
		end
	end
	else
	begin: single_sp_ram_gen
`ifdef FPGA_SRAM
`ifdef ALTERA_EP4
		altera_sp_sram_gen
		#(
			.ADDR_WIDTH(ADDR_WIDTH),
			.DATA_WIDTH(FULL_DATA_WIDTH),
			.BYTE_WIDTH(BYTE_WIDTH),
			.MEM_INITFILE(),
			.DEVICE_FAMILY("Cyclone IV E")
		)
		u_sp_sram_gen
		(
			.clk						(clk),
			.rst						(rst),
			.byteena					(be),
			.wren						(we&cs),
			.rden						(!we&cs)),//?
			.addr						(addr),
			.data						(real_data),
			.q							(real_q)
		);
`elsif ZYNQ_7020
		xilinx_sp_sram_gen
		#(
			.ADDR_WIDTH(ADDR_WIDTH),
			.DATA_WIDTH(FULL_DATA_WIDTH),
			.BYTE_WIDTH(BYTE_WIDTH),
			.MEM_INITFILE(),
			.DEVICE_FAMILY("ZYNQ_7020")
		)
		u_sp_sram_gen
		(
			.clk						(clk),
			.rst						(rst),
			.wea						({BYTE_NUMBER{we}}&be),
			.ena						(cs),
			.addr						(addr),
			.data						(real_data),
			.q							(real_q)
		);
`else
`endif
`else
		sim_sp_sram_gen
		#(
			.ADDR_WIDTH(ADDR_WIDTH),
			.DATA_WIDTH(FULL_DATA_WIDTH),
			.BYTE_WIDTH(BYTE_WIDTH),
			.MEM_INITFILE(),
			.DEVICE_FAMILY("ZYNQ_7020")
		)
		u_sp_sram_gen
		(
			.clk						(clk),
			.rst						(rst),
			.wea						({BYTE_NUMBER{we}}&be),
			.ena						(cs),
			.addr						(addr),
			.data						(real_data),
			.q							(real_q)
		);
`endif
	end
endgenerate


endmodule

