//===============================================
//
//	File: mcu_top.v
//	Author: afterGlow,4ever
//	Group: Fall For Laboratory
//	Date: 07022023
//	Version: v1.0
//
// 	This is top for mcu 'cm3_ahbmtx'.
//	This top is including:
//	ao domain: Always on domain.
//	fp domain: Full function domain.
//	pad top: Ports top.
//	fpga top: Only used in fpga platform.
//
//===============================================

module mcu_top 
(
	// debug port group
	input  wire						CLK,  
	input  wire						RSTN,
	input  wire						TDI, 
	input  wire						TCK, 
	inout  wire						TMS, 
	output wire						TDO, 
	input  wire						TRST 
);

//===============================================
// Top for full function domain
//===============================================
fp_domain u_fp_domain
(
	.sys_root_clk					(CLK				),
	.sys_root_rstn				(RSTN				),
	.apb1_root_clk				(CLK				),
	.apb1_root_rstn				(RSTN				),
	.power_on_rstn				(RSTN				),

	.TDI									(TDI				),
	.TCK									(TCK				),
	.TMS									(TMS				),
	.TDO									(TDO				),
	.TRST									(TRST				)
);

endmodule

