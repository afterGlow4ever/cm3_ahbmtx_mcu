//===============================================
//
//	File: apb2_top.v
//	Author: afterGlow,4ever
//	Group: Fall For Laboratory
//	Date: 02272024
//	Version: v1.0
//
// 	This is top for apb2 async peripherals domain.
//	This domain is including:
//	1. ethernet
//	2. advtim
//	3. spi master
//
//===============================================

module apb2_top 
(
	input						apb2_root_clk,
	input						apb2_root_rstn,
	input  						eth_pe_tx_clk,  
	input  						eth_pe_tx_rstn,
	input  						eth_pe_rx_clk,  
	input  						eth_pe_rx_rstn,
	input  						advtim_pe_clk,  
	input  						advtim_pe_rstn,
	input  						spim_pe_clk,  
	input  						spim_pe_rstn,
	
	// pin
	output 						eth_mdc,
	output 						eth_mdc_oen,
	output 						eth_mdio_o,
	input 						eth_mdio_i,
	output 						eth_mdio_oen,
	output 		[ 3:0]			eth_tx,
	output 		[ 3:0]			eth_tx_oen,
	output 						eth_tx_ctrl,
	output 						eth_tx_ctrl_oen,
	output						eth_tx_clk,	
	output						eth_tx_clk_oen,	
	output						advtmr0_pwm_ch1p,
	output						advtmr0_pwm_ch1n,
	output						advtmr0_pwm_ch2p,
	output						advtmr0_pwm_ch2n,
	output						advtmr0_pwm_ch3p,
	output						advtmr0_pwm_ch3n,
	output						advtmr0_pwm_ch4,
	output						advtmr0_pwm_ch5,
	output						advtmr0_pwm_ch6,
	output						advtmr0_pwm_ch1p_oen,
	output						advtmr0_pwm_ch1n_oen,
	output						advtmr0_pwm_ch2p_oen,
	output						advtmr0_pwm_ch2n_oen,
	output						advtmr0_pwm_ch3p_oen,
	output						advtmr0_pwm_ch3n_oen,
	output						advtmr0_pwm_ch4_oen,
	output						advtmr0_pwm_ch5_oen,
	output						advtmr0_pwm_ch6_oen,
	input						advtmr0_bk1,
	input						advtmr0_bk2,
	output						advtmr0_bk1_oen,
	output						advtmr0_bk2_oen,
	input						advtmr0_cap_ch1p,
	input						advtmr0_cap_ch1n,
	output						advtmr0_cap_ch1p_oen,
	output						advtmr0_cap_ch1n_oen,
	input						advtmr0_enc_ch1p,
	input						advtmr0_enc_ch1n,
	output						advtmr0_enc_ch1p_oen,
	output						advtmr0_enc_ch1n_oen,
	output 						spim0_sck,
	output 						spim0_sck_oen,
	output 						spim0_mosi_o,
	output 						spim0_mosi_oen,
	input						spim0_miso_i,
	output 						spim0_miso_oen,
	output 						spim0_cs_o,
	output 						spim0_cs_oen,

	// event
	input						system_failure,

	// ahb bus
	input						eth_hclk,
	input						eth_hrstn,
	output						eth_hsel,
	output						eth_hreadyout,
	output	[ 1:0]				eth_htrans,
	output	[ 2:0]				eth_hsize,
	output						eth_hwrite,
	output	[ 2:0]				eth_hburst,
	output	[31:0]				eth_haddr,
	output	[ 3:0]				eth_hprot,
	output	[31:0]				eth_hwdata,
	input						eth_hready,
	input	[ 1:0]				eth_hresp,
	input	[31:0]				eth_hrdata,	

	// apb bus
	input	[31:0]				paddr,  
	input						penable,
	input	[ 3:0]				pstrb,  
	input	[ 2:0]				pprot,  
	input						pwrite, 
	input	[31:0]				pwdata, 
	input						psel,   
	output	[31:0]				prdata, 
	output						pready,
	output						pslverr,

	// interrupt line
	output						eth_sma_int,
	output						eth_mac_tx_int,
	output						eth_mac_rx_int,
	output						eth_mac_dma_int,
	output						advtim0_gen_int,
	output						advtim0_cap_int,
	output						advtim0_enc_int,
	output						spim0_int
);

//===============================================
// APB2 slave mux
//===============================================

wire						 	psel_eth; 
wire						 	pready_eth; 
wire	[31:0]				 	prdata_eth; 
wire						 	pslverr_eth; 
wire	[31:0]				 	paddr_eth; 
wire						 	psel_advtim; 
wire						 	pready_advtim; 
wire	[31:0]				 	prdata_advtim; 
wire						 	pslverr_advtim; 
wire	[31:0]				 	paddr_advtim; 
wire						 	psel_spim; 
wire						 	pready_spim; 
wire	[31:0]				 	prdata_spim; 
wire						 	pslverr_spim; 
wire	[31:0]				 	paddr_spim; 

cmsdk_apb_slave_mux 
#(
    .PORT0_ENABLE                       (1),
    .PORT1_ENABLE                       (1),
    .PORT2_ENABLE                       (1),
    .PORT3_ENABLE                       (0),
    .PORT4_ENABLE                       (0),
    .PORT5_ENABLE                       (0),
    .PORT6_ENABLE                       (0),
    .PORT7_ENABLE                       (0),
    .PORT8_ENABLE                       (0),
    .PORT9_ENABLE                       (0),
    .PORT10_ENABLE                      (0),
    .PORT11_ENABLE                      (0),
    .PORT12_ENABLE                      (0),
    .PORT13_ENABLE                      (0),
    .PORT14_ENABLE                      (0),
    .PORT15_ENABLE                      (0)
)   
u_apb2_slave_mux
(
    .DECODE4BIT                         (paddr[15:12]),
    .PSEL                               (psel),

    .PSEL0                              (psel_eth),
    .PREADY0                            (pready_eth),
    .PRDATA0                            (prdata_eth),
    .PSLVERR0                           (pslverr_eth),
    
    .PSEL1                              (psel_advtim),
    .PREADY1                            (pready_advtim),
    .PRDATA1                            (prdata_advtim),
    .PSLVERR1                           (pslverr_advtim),

    .PSEL2                              (psel_spim),
    .PREADY2                            (pready_spim),
    .PRDATA2                            (prdata_spim),
    .PSLVERR2                           (pslverr_spim),

    .PSEL3                              (),
    .PREADY3                            (1'b0),
    .PRDATA3                            (32'b0),
    .PSLVERR3                           (1'b0),

    .PSEL4                              (),
    .PREADY4                            (1'b0),
    .PRDATA4                            (32'b0),
    .PSLVERR4                           (1'b0),

    .PSEL5                              (),
    .PREADY5                            (1'b0),
    .PRDATA5                            (32'b0),
    .PSLVERR5                           (1'b0),

    .PSEL6                              (),
    .PREADY6                            (1'b0),
    .PRDATA6                            (32'b0),
    .PSLVERR6                           (1'b0),

    .PSEL7                              (),
    .PREADY7                            (1'b0),
    .PRDATA7                            (32'b0),
    .PSLVERR7                           (1'b0),

    .PSEL8                              (),
    .PREADY8                            (1'b0),
    .PRDATA8                            (32'b0),
    .PSLVERR8                           (1'b0),

    .PSEL9                              (),
    .PREADY9                            (1'b0),
    .PRDATA9                            (32'b0),
    .PSLVERR9                           (1'b0),

    .PSEL10                             (),
    .PREADY10                           (1'b0),
    .PRDATA10                           (32'b0),
    .PSLVERR10                          (1'b0),

    .PSEL11                             (),
    .PREADY11                           (1'b0),
    .PRDATA11                           (32'b0),
    .PSLVERR11                          (1'b0),

    .PSEL12                             (),
    .PREADY12                           (1'b0),
    .PRDATA12                           (32'b0),
    .PSLVERR12                          (1'b0),
    
    .PSEL13                             (),
    .PREADY13                           (1'b0),
    .PRDATA13                           (32'b0),
    .PSLVERR13                          (1'b0),

    .PSEL14                             (),
    .PREADY14                           (1'b0),
    .PRDATA14                           (32'b0),
    .PSLVERR14                          (1'b0),

    .PSEL15                             (),
    .PREADY15                           (1'b0),
    .PRDATA15                           (32'b0),
    .PSLVERR15                          (1'b0),

    .PREADY                             (pready),
    .PRDATA                             (prdata),
    .PSLVERR                            (pslverr)

);

//===============================================
// APB2 ethernet
// 0x40020000~0x40020FFF 
//===============================================

assign pready_eth = 1'b1;
assign pslverr_eth = 1'b0;

`ifdef ETH
assign paddr_eth = paddr;// compatible with ethernet reg

eth_top u_eth
(
	.module_clk					(apb2_root_clk),  
	.module_rstn				(apb2_root_rstn),
	.pe_tx_clk					(eth_pe_tx_clk),  
	.pe_tx_rstn					(eth_pe_tx_rstn),
	.pe_rx_clk					(eth_pe_rx_clk),  
	.pe_rx_rstn					(eth_pe_rx_rstn),

	.eth_mdc					(eth_mdc),
	.eth_mdc_oen				(eth_mdc_oen),
	.eth_mdio_o					(eth_mdio_o),
	.eth_mdio_i					(eth_mdio_i),
	.eth_mdio_oen				(eth_mdio_oen),
	.eth_tx						(eth_tx),
	.eth_tx_oen					(eth_tx_oen),
	.eth_tx_ctrl				(eth_tx_ctrl),
	.eth_tx_ctrl_oen			(eth_tx_ctrl_oen),
	.eth_tx_clk					(eth_tx_clk),	
	.eth_tx_clk_oen				(eth_tx_clk_oen),	

	.ahb_hclk					(eth_hclk),
	.ahb_hrstn					(eth_hrstn),
	.ahb_hsel					(eth_hsel),
	.ahb_hreadyout				(eth_hreadyout),
	.ahb_htrans					(eth_htrans),
	.ahb_hsize					(eth_hsize),
	.ahb_hwrite					(eth_hwrite),
	.ahb_hburst					(eth_hburst),
	.ahb_haddr					(eth_haddr),
	.ahb_hprot					(eth_hprot),
	.ahb_hwdata					(eth_hwdata),
	.ahb_hready					(eth_hready),
	.ahb_hresp					(eth_hresp),
	.ahb_hrdata					(eth_hrdata),	

	.reg_clk					(apb2_root_clk),
	.reg_rstn					(apb2_root_rstn),
	.pwrite						(pwrite),
	.psel						(psel_eth),						
	.penable					(penable),
	.paddr						(paddr_eth),
	.pwdata						(pwdata),
	.prdata						(prdata_eth),

	.eth_sma_int_line			(eth_sma_int),
	.eth_mac_tx_int_line		(eth_mac_tx_int),
	.eth_mac_rx_int_line		(eth_mac_rx_int),
	.eth_mac_dma_int_line		(eth_mac_dma_int)
);
`else
assign eth_mdc = 1'b0;
assign eth_mdc_oen = 1'b0;
assign eth_mdio_o = 1'b0;
assign eth_mdio_oen = 1'b0;
assign eth_tx = 4'h0;
assign eth_tx_oen = 4'h0;
assign eth_tx_ctrl = 1'b0;	
assign eth_tx_ctrl_oen = 1'b0;
assign eth_tx_clk = 1'b0;		
assign eth_tx_clk_oen = 1'b0;	
assign eth_haddr = 32'h0;
assign eth_htrans = 2'h0;
assign eth_hsize = 3'h0;
assign eth_hwrite = 1'b0;
assign eth_hwdata = 32'h0;
assign eth_hreadyout = 1'b1;
assign prdata_eth = 32'h0;
assign eth_sma_int = 1'b0;
assign eth_mac_tx_int = 1'b0;
assign eth_mac_rx_int = 1'b0;
assign eth_mac_dma_int = 1'b0;
`endif

//===============================================
// APB2 advance timer
// 0x40021000~0x40021FFF 
//===============================================

assign pready_advtim = 1'b1;
assign pslverr_advtim = 1'b0;

`ifdef ADVTIM
assign paddr_advtim = paddr;// compatible with advanve timer reg

advtim_top u_advtim
(
	.module_clk					(advtim_pe_clk),  
	.module_rstn				(advtim_pe_rstn),

	.advtmr_pwm_ch1p			(advtmr0_pwm_ch1p),
	.advtmr_pwm_ch1n			(advtmr0_pwm_ch1n),
	.advtmr_pwm_ch2p			(advtmr0_pwm_ch2p),
	.advtmr_pwm_ch2n			(advtmr0_pwm_ch2n),
	.advtmr_pwm_ch3p			(advtmr0_pwm_ch3p),
	.advtmr_pwm_ch3n			(advtmr0_pwm_ch3n),
	.advtmr_pwm_ch4				(advtmr0_pwm_ch4),
	.advtmr_pwm_ch5				(advtmr0_pwm_ch5),
	.advtmr_pwm_ch6				(advtmr0_pwm_ch6),
	.advtmr_pwm_ch1p_oen		(advtmr0_pwm_ch1p_oen),
	.advtmr_pwm_ch1n_oen		(advtmr0_pwm_ch1n_oen),
	.advtmr_pwm_ch2p_oen		(advtmr0_pwm_ch2p_oen),
	.advtmr_pwm_ch2n_oen		(advtmr0_pwm_ch2n_oen),
	.advtmr_pwm_ch3p_oen		(advtmr0_pwm_ch3p_oen),
	.advtmr_pwm_ch3n_oen		(advtmr0_pwm_ch3n_oen),
	.advtmr_pwm_ch4_oen			(advtmr0_pwm_ch4_oen),
	.advtmr_pwm_ch5_oen			(advtmr0_pwm_ch5_oen),
	.advtmr_pwm_ch6_oen			(advtmr0_pwm_ch6_oen),
	.advtmr_bk1					(advtmr0_bk1),
	.advtmr_bk2					(advtmr0_bk2),
	.advtmr_bk1_oen				(advtmr0_bk1_oen),
	.advtmr_bk2_oen				(advtmr0_bk2_oen),
	.advtmr_cap_ch1p			(advtmr0_cap_ch1p),
	.advtmr_cap_ch1n			(advtmr0_cap_ch1n),
	.advtmr_cap_ch1p_oen		(advtmr0_cap_ch1p_oen),
	.advtmr_cap_ch1n_oen		(advtmr0_cap_ch1n_oen),
	.advtmr_enc_ch1p			(advtmr0_enc_ch1p),
	.advtmr_enc_ch1n			(advtmr0_enc_ch1n),
	.advtmr_enc_ch1p_oen		(advtmr0_enc_ch1p_oen),
	.advtmr_enc_ch1n_oen		(advtmr0_enc_ch1n_oen),

	.system_failure				(system_failure),

	.reg_clk					(apb2_root_clk),
	.reg_rstn					(apb2_root_rstn),
	.pwrite						(pwrite),
	.psel						(psel_advtim),						
	.penable					(penable),
	.paddr						(paddr_advtim),
	.pwdata						(pwdata),
	.prdata						(prdata_advtim),

	.advtim_gen_int_line		(advtim0_gen_int),
	.advtim_cap_int_line		(advtim0_cap_int),
	.advtim_enc_int_line		(advtim0_enc_int)
);
`else
assign advtmr0_pwm_ch1p = 1'b0;
assign advtmr0_pwm_ch1n = 1'b0;
assign advtmr0_pwm_ch2p = 1'b0;
assign advtmr0_pwm_ch2n = 1'b0;
assign advtmr0_pwm_ch3p = 1'b0;
assign advtmr0_pwm_ch3n = 1'b0;
assign advtmr0_pwm_ch4 = 1'b0;
assign advtmr0_pwm_ch5 = 1'b0;
assign advtmr0_pwm_ch6 = 1'b0;
assign advtmr0_pwm_ch1p_oen = 1'b0;
assign advtmr0_pwm_ch1n_oen = 1'b0;
assign advtmr0_pwm_ch2p_oen = 1'b0;
assign advtmr0_pwm_ch2n_oen = 1'b0;
assign advtmr0_pwm_ch3p_oen = 1'b0;
assign advtmr0_pwm_ch3n_oen = 1'b0;
assign advtmr0_pwm_ch4_oen = 1'b0;
assign advtmr0_pwm_ch5_oen = 1'b0;
assign advtmr0_pwm_ch6_oen = 1'b0;
assign advtmr0_bk1_oen = 1'b0;
assign advtmr0_bk2_oen = 1'b0;
assign advtmr0_cap_ch1p_oen = 1'b0;
assign advtmr0_cap_ch1n_oen = 1'b0;
assign prdata_advtim = 32'h0;
assign advtim0_gen_int = 1'b0;
assign advtim0_cap_int = 1'b0;
assign advtim0_enc_int = 1'b0;
`endif

//===============================================
// APB2 spi master
// 0x40022000~0x40022FFF
//===============================================

assign pready_spim = 1'b1;
assign pslverr_spim = 1'b0;

`ifdef SPIM
assign paddr_spim = paddr;// compatible with uart reg

spim_top u_spim
(
	.module_clk					(spim_pe_clk),  
	.module_rstn				(spim_pe_rstn),
	
	.spim_sck					(spim0_sck),
	.spim_sck_oen				(spim0_sck_oen),
	.spim_mosi_o				(spim0_mosi_o),
	.spim_mosi_oen				(spim0_mosi_oen),
	.spim_miso_i				(spim0_miso_i),
	.spim_miso_oen				(spim0_miso_oen),
	.spim_cs_o					(spim0_cs_o),
	.spim_cs_oen				(spim0_cs_oen),

	.reg_clk					(apb2_root_clk),
	.reg_rstn					(apb2_root_rstn),
	.pwrite						(pwrite),
	.psel						(psel_spim),						
	.penable					(penable),
	.paddr						(paddr_spim),
	.pwdata						(pwdata),
	.prdata						(prdata_spim),

	.spim_int_line				(spim0_int)
);
`else
assign spim0_sck = 1'b0;
assign spim0_sck_oen = 1'b0;
assign spim0_mosi_o = 1'b0;
assign spim0_mosi_oen = 1'b0;
assign prdata_spim = 32'h0;
assign spim0_int = 1'b0;
`endif


endmodule

